--not R0, R1