--div R6, R7