--OR R1, R2, R3