--add R0, R4, R5