--shr R1, R3, R5