--mul R6, R7