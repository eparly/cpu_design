--neg R0, R1