--ror R6, R6, R4